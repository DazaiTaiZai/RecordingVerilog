module latches (

);
    
endmodule